`timescale 1 ns / 1 ps
//
`default_nettype none

module rs_encoder (
    input  wire       clk,
    input  wire       rst_n,
    //
    input  wire [7:0] msg_in      [64],
    input  wire       msg_valid,
    //
    output wire [7:0] parity_out  [ 4],
    output wire       parity_valid
);

  // verilog_format: off
  logic [7:0] log_table [256] = '{
     -1,   0,   1,  25,   2,  50,  26, 198,   3, 223,  51, 238,  27, 104, 199,  75,
      4, 100, 224,  14,  52, 141, 239, 129,  28, 193, 105, 248, 200,   8,  76, 113,
      5, 138, 101,  47, 225,  36,  15,  33,  53, 147, 142, 218, 240,  18, 130,  69,
     29, 181, 194, 125, 106,  39, 249, 185, 201, 154,   9, 120,  77, 228, 114, 166,
      6, 191, 139,  98, 102, 221,  48, 253, 226, 152,  37, 179,  16, 145,  34, 136,
     54, 208, 148, 206, 143, 150, 219, 189, 241, 210,  19,  92, 131,  56,  70,  64,
     30,  66, 182, 163, 195,  72, 126, 110, 107,  58,  40,  84, 250, 133, 186,  61,
    202,  94, 155, 159,  10,  21, 121,  43,  78, 212, 229, 172, 115, 243, 167,  87,
      7, 112, 192, 247, 140, 128,  99,  13, 103,  74, 222, 237,  49, 197, 254,  24,
    227, 165, 153, 119,  38, 184, 180, 124,  17,  68, 146, 217,  35,  32, 137,  46,
     55,  63, 209,  91, 149, 188, 207, 205, 144, 135, 151, 178, 220, 252, 190,  97,
    242,  86, 211, 171,  20,  42,  93, 158, 132,  60,  57,  83,  71, 109,  65, 162,
     31,  45,  67, 216, 183, 123, 164, 118, 196,  23,  73, 236, 127,  12, 111, 246,
    108, 161,  59,  82,  41, 157,  85, 170, 251,  96, 134, 177, 187, 204,  62,  90,
    203,  89,  95, 176, 156, 169, 160,  81,  11, 245,  22, 235, 122, 117,  44, 215,
     79, 174, 213, 233, 230, 231, 173, 232, 116, 214, 244, 234, 168,  80,  88, 175
  };

  reg [7:0] exp_table [256] = '{
      1,   2,   4,   8,  16,  32,  64, 128,  29,  58, 116, 232, 205, 135,  19,  38,
     76, 152,  45,  90, 180, 117, 234, 201, 143,   3,   6,  12,  24,  48,  96, 192,
    157,  39,  78, 156,  37,  74, 148,  53, 106, 212, 181, 119, 238, 193, 159,  35,
     70, 140,   5,  10,  20,  40,  80, 160,  93, 186, 105, 210, 185, 111, 222, 161,
     95, 190,  97, 194, 153,  47,  94, 188, 101, 202, 137,  15,  30,  60, 120, 240,
    253, 231, 211, 187, 107, 214, 177, 127, 254, 225, 223, 163,  91, 182, 113, 226,
    217, 175,  67, 134,  17,  34,  68, 136,  13,  26,  52, 104, 208, 189, 103, 206,
    129,  31,  62, 124, 248, 237, 199, 147,  59, 118, 236, 197, 151,  51, 102, 204,
    133,  23,  46,  92, 184, 109, 218, 169,  79, 158,  33,  66, 132,  21,  42,  84,
    168,  77, 154,  41,  82, 164,  85, 170,  73, 146,  57, 114, 228, 213, 183, 115,
    230, 209, 191,  99, 198, 145,  63, 126, 252, 229, 215, 179, 123, 246, 241, 255,
    227, 219, 171,  75, 150,  49,  98, 196, 149,  55, 110, 220, 165,  87, 174,  65,
    130,  25,  50, 100, 200, 141,   7,  14,  28,  56, 112, 224, 221, 167,  83, 166,
     81, 162,  89, 178, 121, 242, 249, 239, 195, 155,  43,  86, 172,  69, 138,   9,
     18,  36,  72, 144,  61, 122, 244, 245, 247, 243, 251, 235, 203, 139,  11,  22,
     44,  88, 176, 125, 250, 233, 207, 131,  27,  54, 108, 216, 173,  71, 142,  -1
  };

  reg [7:0] g_table [64][4] = '{
    {174,  27, 162,  37},
    { 27, 212, 123,  61},
    { 51,  31,  19, 243},
    {233,  19,  57, 103},
    { 93, 239,  83, 179},
    {169,  64,  13, 170},
    {160, 130,  83,  90},
    { 80,   1,  29,  40},
    { 30,  23,   2,  88},
    { 78, 210,   6,  43},
    { 33, 123,  58, 167},
    {157,  41, 189, 182},
    {172, 111,  53,   4},
    {249,  36,  33,  33},
    { 23, 242,  87, 142},
    {132,  17,  39, 197},
    {187, 188, 131, 211},
    {201, 249,  53,  54},
    { 44,  25, 131, 248},
    {238,  77, 116,  25},
    { 15, 144,  41, 138},
    {128, 234, 166, 121},
    {111, 210, 119, 109},
    { 99, 181,  83,  50},
    { 40, 167,  52,  12},
    {  2, 224, 154,  97},
    { 87, 110, 135, 123},
    {113,  53, 134, 217},
    {207, 198, 196,  80},
    { 70,  77, 126, 182},
    {172, 221,  31, 138},
    {128, 207,  59, 182},
    {172, 137,  19, 184},
    {174, 129, 152,  92},
    { 82,  48,  61, 142},
    {132, 192, 216,  32},
    { 22, 234,  97, 179},
    {169,  25,  40, 216},
    {206, 245, 159, 232},
    {222, 225,  67,  39},
    { 29, 227,  33, 188},
    {178,  65,  66, 185},
    {175, 159, 104, 163},
    {153, 128, 170, 173},
    {163, 140, 173,  18},
    {  8,   3,  38, 129},
    {119, 212,  10, 103},
    { 93, 121,  17, 128},
    {118, 140, 226, 180},
    {170,   3,  83, 227},
    {217,  98, 244, 127},
    {117, 192, 131,  80},
    { 70,  43, 176, 173},
    {163, 226,   2, 193},
    {183, 159,  25, 114},
    {104, 148, 182, 106},
    { 96, 121, 223,  60},
    { 50, 162, 245, 150},
    {140, 164,  79, 220},
    {210, 102, 184, 157},
    {147,  54,   4, 144},
    {134, 202, 167, 175},
    {165, 192,  63,  86},
    { 76, 251,  81,  10}
  };
  // verilog_format: on


  logic [7:0] log_msg[64];
  logic       msg_z  [64];

  logic [8:0] mul0[64][4];
  logic [7:0] mul1[64][4];
  logic [7:0] mul2[64][4];

  logic [7:0] add   [4];
  logic [7:0] parity[4];
  logic       valid;

  generate
    for (genvar i = 0; i < 64; i++) begin

      assign log_msg[i] = log_table[msg_in[i]];
      assign msg_z[i]   = (msg_in[i] == 0);

      for (genvar j = 0; j < 4; j++) begin

        assign mul0[i][j] = log_msg[i] + g_table[i][j];

        assign mul1[i][j] = (mul0[i][j] >= 255) ? (mul0[i][j] - 255) : mul0[i][j];

        assign mul2[i][j] = msg_z[i] ? '0 : exp_table[mul1[i][j]];

      end

    end
  endgenerate

  generate
    for (genvar j = 0; j < 4; j++) begin

      always_comb begin
        add[j] = '0;
        for (int i = 0; i < 64; i++) begin
          add[j] = add[j] ^ mul2[i][j];
        end
      end

      always_ff @(posedge clk) begin
        parity[j] <= add[j];
      end

      assign parity_out[j] = parity[j];

    end
  endgenerate

  always_ff @(posedge clk) begin
    valid <= msg_valid;
  end

  assign parity_valid = valid;

endmodule

`default_nettype wire
