`timescale 1 ns / 1 ps
//
`default_nettype none

module rs_encoder (
    input  wire       clk,
    input  wire       rst_n,
    //
    input  wire [7:0] msg_in    [64],
    input  wire       vld_in,
    //
    output wire [7:0] msg_out   [64],
    output wire [7:0] parity_out[ 4],
    output wire       vld_out
);

  localparam logic [7:0] prim = 8'h1d;

  // verilog_format: off
  localparam logic [7:0] g_table_a0 [64][4] = '{
    {241,  12, 191,  74},
    { 12, 121, 197, 111},
    { 10, 192,  90, 125},
    {243,  90, 186, 136},
    {182,  22, 187,  75},
    {229,  95, 135, 215},
    {230,  46, 187, 223},
    {253,   2,  48, 106},
    { 96, 201,   4, 254},
    {120,  89,  64, 119},
    { 39, 197, 105, 126},
    {213, 212,  87,  98},
    {123, 206,  40,  16},
    { 54,  37,  39,  39},
    {201, 176, 127,  42},
    {184, 152,  53, 141},
    {220, 165,  92, 178},
    { 56,  54,  40,  80},
    {238,   3,  92,  27},
    { 11,  60, 248,   3},
    { 38, 168, 212,  33},
    {133, 251,  63, 118},
    {206,  89, 147, 189},
    {134,  49, 187,   5},
    {106, 126,  20, 205},
    {  4,  18,  57, 175},
    {127, 103, 169, 197},
    { 31,  40, 218, 155},
    {166,   7, 200, 253},
    { 94,  60, 102,  98},
    {123,  69, 192,  33},
    {133, 166, 210,  98},
    {123, 158,  90, 149},
    {241,  23,  73,  91},
    {211,  70, 111,  42},
    {184, 130, 195, 157},
    {234, 251, 175,  75},
    {229,   3, 106, 195},
    { 83, 233, 115, 247},
    {138,  36, 194,  53},
    { 48, 144,  39, 165},
    {171, 190,  97,  55},
    {255, 115,  13,  99},
    {146, 133, 215, 246},
    { 99, 132, 246,  45},
    { 29,   8, 148,  23},
    {147, 121, 116, 136},
    {182, 118, 152, 133},
    {199, 132,  72, 150},
    {215,   8, 187, 144},
    {155,  67, 250, 204},
    {237, 130,  92, 253},
    { 94, 119, 227, 246},
    { 99,  72,   4,  25},
    {196, 115,   3,  62},
    { 13,  82,  98,  52},
    {217, 118,   9, 185},
    {  5, 191, 233,  85},
    {132, 198, 240, 172},
    { 89,  68, 149, 213},
    { 41,  80,  16, 168},
    {218, 112, 126, 255},
    {145, 130, 161, 177},
    { 30, 216, 231, 116}
  };

  localparam logic [7:0] g_table_a1 [64][4] = '{
    {255,  24,  99, 148},
    { 24, 242, 151, 222},
    { 20, 157, 180, 250},
    {251, 180, 105,  13},
    {113,  44, 107, 150},
    {215, 190,  19, 179},
    {209,  92, 107, 163},
    {231,   4,  96, 212},
    {192, 143,   8, 225},
    {240, 178, 128, 238},
    { 78, 151, 210, 252},
    {183, 181, 174, 196},
    {246, 129,  80,  32},
    {108,  74,  78,  78},
    {143, 125, 254,  84},
    {109,  45, 106,   7},
    {165,  87, 184, 121},
    {112, 108,  80, 160},
    {193,   6, 184,  54},
    { 22, 120, 237,   6},
    { 76,  77, 181,  66},
    { 23, 235, 126, 236},
    {129, 178,  59, 103},
    { 17,  98, 107,  10},
    {212, 252,  40, 135},
    {  8,  36, 114,  67},
    {254, 206,  79, 151},
    { 62,  80, 169,  43},
    { 81,  14, 141, 231},
    {188, 120, 204, 196},
    {246, 138, 157,  66},
    { 23,  81, 185, 196},
    {246,  33, 180,  55},
    {255,  46, 146, 182},
    {187, 140, 222,  84},
    {109,  25, 155,  39},
    {201, 235,  67, 150},
    {215,   6, 212, 155},
    {166, 207, 230, 243},
    {  9,  72, 153, 106},
    { 96,  61,  78,  87},
    { 75,  97, 194, 110},
    {227, 230,  26, 198},
    { 57,  23, 179, 241},
    {198,  21, 241,  90},
    { 58,  16,  53,  46},
    { 59, 242, 232,  13},
    {113, 236,  45,  23},
    {147,  21, 144,  49},
    {179,  16, 107,  61},
    { 43, 134, 233, 133},
    {199,  25, 184, 231},
    {188, 238, 219, 241},
    {198, 144,   8,  50},
    {149, 230,   6, 124},
    { 26, 164, 196, 104},
    {175, 236,  18, 111},
    { 10,  99, 207, 170},
    { 21, 145, 253,  69},
    {178, 136,  55, 183},
    { 82, 160,  32,  77},
    {169, 224, 252, 227},
    { 63,  25,  95, 127},
    { 60, 173, 211, 232}
  };

  localparam logic [7:0] g_table_a2 [64][4] = '{
    {227,  48, 198,  53},
    { 48, 249,  51, 161},
    { 40,  39, 117, 233},
    {235, 117, 210,  26},
    {226,  88, 214,  49},
    {179,  97,  38, 123},
    {191, 184, 214,  91},
    {211,   8, 192, 181},
    {157,   3,  16, 223},
    {253, 121,  29, 193},
    {156,  51, 185, 229},
    {115, 119,  65, 149},
    {241,  31, 160,  64},
    {216, 148, 156, 156},
    {  3, 250, 225, 168},
    {218,  90, 212,  14},
    { 87, 174, 109, 242},
    {224, 216, 160,  93},
    {159,  12, 109, 108},
    { 44, 240, 199,  12},
    {152, 154, 119, 132},
    { 46, 203, 252, 197},
    { 31, 121, 118, 206},
    { 34, 196, 214,  20},
    {181, 229,  80,  19},
    { 16,  72, 228, 134},
    {225, 129, 158,  51},
    {124, 160,  79,  86},
    {162,  28,   7, 211},
    {101, 240, 133, 149},
    {241,   9,  39, 132},
    { 46, 162, 111, 149},
    {241,  66, 117, 110},
    {227,  92,  57, 113},
    {107,   5, 161, 168},
    {218,  50,  43,  78},
    {143, 203, 134,  49},
    {179,  12, 181,  43},
    { 81, 131, 209, 251},
    { 18, 144,  47, 212},
    {192, 122, 156, 174},
    {150, 194, 153, 220},
    {219, 209,  52, 145},
    {114,  46, 123, 255},
    {145,  42, 255, 180},
    {116,  32, 106,  92},
    {118, 249, 205,  26},
    {226, 197,  90,  46},
    { 59,  42,  61,  98},
    {123,  32, 214, 122},
    { 86,  17, 207,  23},
    {147,  50, 109, 211},
    {101, 193, 171, 255},
    {145,  61,  16, 100},
    { 55, 209,  12, 248},
    { 52,  85, 149, 208},
    { 67, 197,  36, 222},
    { 20, 198, 131,  73},
    { 42,  63, 231, 138},
    {121,  13, 110, 115},
    {164,  93,  64, 154},
    { 79, 221, 229, 219},
    {126,  50, 190, 254},
    {120,  71, 187, 205}
  };

  localparam logic [7:0] g_table_a3 [64][4] = '{
    {219,  96, 145, 106},
    { 96, 239, 102,  95},
    { 80,  78, 234, 207},
    {203, 234, 185,  52},
    {217, 176, 177,  98},
    {123, 194,  76, 246},
    { 99, 109, 177, 182},
    {187,  16, 157, 119},
    { 39,   6,  32, 163},
    {231, 242,  58, 159},
    { 37, 102, 111, 215},
    {230, 238, 130,  55},
    {255,  62,  93, 128},
    {173,  53,  37,  37},
    {  6, 233, 223,  77},
    {169, 180, 181,  28},
    {174,  65, 218, 249},
    {221, 173,  93, 186},
    { 35,  24, 218, 216},
    { 88, 253, 147,  24},
    { 45,  41, 238,  21},
    { 92, 139, 229, 151},
    { 62, 242, 236, 129},
    { 68, 149, 177,  40},
    {119, 215, 160,  38},
    { 32, 144, 213,  17},
    {223,  31,  33, 102},
    {248,  93, 158, 172},
    { 89,  56,  14, 187},
    {202, 253,  23,  55},
    {255,  18,  78,  21},
    { 92,  89, 222,  55},
    {255, 132, 234, 220},
    {219, 184, 114, 226},
    {214,  10,  95,  77},
    {169, 100,  86, 156},
    {  3, 139,  17,  98},
    {123,  24, 119,  86},
    {162,  27, 191, 235},
    { 36,  61,  94, 181},
    {157, 244,  37,  65},
    { 49, 153,  47, 165},
    {171, 191, 104,  63},
    {228,  92, 246, 227},
    { 63,  84, 227, 117},
    {232,  64, 212, 184},
    {236, 239, 135,  52},
    {217, 151, 180,  92},
    {118,  84, 122, 196},
    {246,  64, 177, 244},
    {172,  34, 131,  46},
    { 59, 100, 218, 187},
    {202, 159,  75, 227},
    { 63, 122,  32, 200},
    {110, 191,  24, 237},
    {104, 170,  55, 189},
    {134, 151,  72, 161},
    { 40, 145,  27, 146},
    { 84, 126, 211,   9},
    {242,  26, 220, 230},
    { 85, 186, 128,  41},
    {158, 167, 215, 171},
    {252, 100,  97, 225},
    {240, 142, 107, 135}
  };

  localparam logic [7:0] g_table_a4 [64][4] = '{
    {171, 192,  63, 212},
    {192, 195, 204, 190},
    {160, 156, 201, 131},
    {139, 201, 111, 104},
    {175, 125, 127, 196},
    {246, 153, 152, 241},
    {198, 218, 127, 113},
    {107,  32,  39, 238},
    { 78,  12,  64,  91},
    {211, 249, 116,  35},
    { 74, 204, 222, 179},
    {209, 193,  25, 110},
    {227, 124, 186,  29},
    { 71, 106,  74,  74},
    { 12, 207, 163, 154},
    { 79, 117, 119,  56},
    { 65, 130, 169, 239},
    {167,  71, 186, 105},
    { 70,  48, 169, 173},
    {176, 231,  59,  48},
    { 90,  82, 193,  42},
    {184,  11, 215,  51},
    {124, 249, 197,  31},
    {136,  55, 127,  80},
    {238, 179,  93,  76},
    { 64,  61, 183,  34},
    {163,  62,  66, 204},
    {237, 186,  33,  69},
    {178, 112,  28, 107},
    {137, 231,  46, 110},
    {227,  36, 156,  42},
    {184, 178, 161, 110},
    {227,  21, 201, 165},
    {171, 109, 228, 217},
    {177,  20, 190, 154},
    { 79, 200, 172,  37},
    {  6,  11,  34, 196},
    {246,  48, 238, 172},
    { 89,  54,  99, 203},
    { 72, 122, 188, 119},
    { 39, 245,  74, 130},
    { 98,  47,  94,  87},
    { 75,  99, 208, 126},
    {213, 184, 241, 219},
    {126, 168, 219, 234},
    {205, 128, 181, 109},
    {197, 195,  19, 104},
    {175,  51, 117, 184},
    {236, 168, 244, 149},
    {241, 128, 127, 245},
    { 69,  68,  27,  92},
    {118, 200, 169, 107},
    {137,  35, 150, 219},
    {126, 244,  64, 141},
    {220,  99,  48, 199},
    {208,  73, 110, 103},
    { 17,  51, 144,  95},
    { 80,  63,  54,  57},
    {168, 252, 187,  18},
    {249,  52, 165, 209},
    {170, 105,  29,  82},
    { 33,  83, 179,  75},
    {229, 200, 194, 223},
    {253,   1, 214,  19}
  };

  localparam logic [7:0] g_table_a5 [64][4] = '{
    { 75, 157, 126, 181},
    {157, 155, 133,  97},
    { 93,  37, 143,  27},
    { 11, 143, 222, 208},
    { 67, 250, 254, 149},
    {241,  47,  45, 255},
    {145, 169, 254, 226},
    {214,  64,  78, 193},
    {156,  24, 128, 182},
    {187, 239, 232,  70},
    {148, 133, 161, 123},
    {191, 159,  50, 220},
    {219, 248, 105,  58},
    {142, 212, 148, 148},
    { 24, 131,  91,  41},
    {158, 234, 238, 112},
    {130,  25,  79, 195},
    { 83, 142, 105, 210},
    {140,  96,  79,  71},
    {125, 211, 118,  96},
    {180, 164, 159,  84},
    {109,  22, 179, 102},
    {248, 239, 151,  62},
    { 13, 110, 254, 160},
    {193, 123, 186, 152},
    {128, 122, 115,  68},
    { 91, 124, 132, 133},
    {199, 105,  66, 138},
    {121, 224,  56, 214},
    { 15, 211,  92, 220},
    {219,  72,  37,  84},
    {109, 121,  95, 220},
    {219,  42, 143,  87},
    { 75, 218, 213, 175},
    {127,  40,  97,  41},
    {158, 141,  69,  74},
    { 12,  22,  68, 149},
    {241,  96, 193,  69},
    {178, 108, 198, 139},
    {144, 244, 101, 238},
    { 78, 247, 148,  25},
    {196,  94, 188, 174},
    {150, 198, 189, 252},
    {183, 109, 255, 171},
    {252,  77, 171, 201},
    {135,  29, 119, 218},
    {151, 155,  38, 208},
    { 67, 102, 234, 109},
    {197,  77, 245,  55},
    {255,  29, 254, 247},
    {138, 136,  54, 184},
    {236, 141,  79, 214},
    { 15,  70,  49, 171},
    {252, 245, 128,   7},
    {165, 198,  96, 147},
    {189, 146, 220, 206},
    { 34, 102,  61, 190},
    {160, 126, 108, 114},
    { 77, 229, 107,  36},
    {239, 104,  87, 191},
    { 73, 210,  58, 164},
    { 66, 166, 123, 150},
    {215, 141, 153, 163},
    {231,   2, 177,  38}
  };

  localparam logic [7:0] g_table_a6 [64][4] = '{
    {150,  39, 252, 119},
    { 39,  43,  23, 194},
    {186,  74,   3,  54},
    { 22,   3, 161, 189},
    {134, 233, 225,  55},
    {255,  94,  90, 227},
    { 63,  79, 225, 217},
    {177, 128, 156, 159},
    { 37,  48,  29, 113},
    {107, 195, 205, 140},
    { 53,  23,  95, 246},
    { 99,  35, 100, 165},
    {171, 237, 210, 116},
    {  1, 181,  53,  53},
    { 48,  27, 182,  82},
    { 33, 201, 193, 224},
    { 25,  50, 158, 155},
    {166,   1, 210, 185},
    {  5, 192, 158, 142},
    {250, 187, 236, 192},
    {117,  85,  35, 168},
    {218,  44, 123, 204},
    {237, 195,  51, 124},
    { 26, 220, 225,  93},
    {159, 246, 105,  45},
    { 29, 244, 230, 136},
    {182, 248,  21,  23},
    {147, 210, 132,   9},
    {242, 221, 112, 177},
    { 30, 187, 184, 165},
    {171, 144,  74, 168},
    {218, 242, 190, 165},
    {171,  84,   3, 174},
    {150, 169, 183,  67},
    {254,  80, 194,  82},
    { 33,   7, 138, 148},
    { 24,  44, 136,  55},
    {255, 192, 159, 138},
    {121, 216, 145,  11},
    { 61, 245, 202, 193},
    {156, 243,  53,  50},
    {149, 188, 101,  65},
    { 49, 145, 103, 229},
    {115, 218, 227,  75},
    {229, 154,  75, 143},
    { 19,  58, 238, 169},
    { 51,  43,  76, 189},
    {134, 204, 201, 218},
    {151, 154, 247, 110},
    {227,  58, 225, 243},
    {  9,  13, 108, 109},
    {197,   7, 158, 177},
    { 30, 140,  98,  75},
    {229, 247,  29,  14},
    { 87, 145, 192,  59},
    {103,  57, 165, 129},
    { 68, 204, 122,  97},
    { 93, 252, 216, 228},
    {154, 215, 214,  72},
    {195, 208, 174,  99},
    {146, 185, 116,  85},
    {132,  81, 246,  49},
    {179,   7,  47,  91},
    {211,   4, 127,  76}
  };

  localparam logic [7:0] g_table_a7 [64][4] = '{
    { 49,  78, 229, 238},
    { 78,  86,  46, 153},
    {105, 148,   6, 108},
    { 44,   6,  95, 103},
    { 17, 207, 223, 110},
    {227, 188, 180, 219},
    {126, 158, 223, 175},
    {127,  29,  37,  35},
    { 74,  96,  58, 226},
    {214, 155, 135,   5},
    {106,  46, 190, 241},
    {198,  70, 200,  87},
    { 75, 199, 185, 232},
    {  2, 119, 106, 106},
    { 96,  54, 113, 164},
    { 66, 143, 159, 221},
    { 50, 100,  33,  43},
    { 81,   2, 185, 111},
    { 10, 157,  33,   1},
    {233, 107, 197, 157},
    {234, 170,  70,  77},
    {169,  88, 246, 133},
    {199, 155, 102, 248},
    { 52, 165, 223, 186},
    { 35, 241, 210,  90},
    { 58, 245, 209,  13},
    {113, 237,  42,  46},
    { 59, 185,  21,  18},
    {249, 167, 224, 127},
    { 60, 107, 109,  87},
    { 75,  61, 148,  77},
    {169, 249,  97,  87},
    { 75, 168,   6,  65},
    { 49,  79, 115, 134},
    {225, 160, 153, 164},
    { 66,  14,   9,  53},
    { 48,  88,  13, 110},
    {227, 157,  35,   9},
    {242, 173,  63,  22},
    {122, 247, 137, 159},
    { 37, 251, 106, 100},
    { 55, 101, 202, 130},
    { 98,  63, 206, 215},
    {230, 169, 219, 150},
    {215,  41, 150,   3},
    { 38, 116, 193,  79},
    {102,  86, 152, 103},
    { 17, 133, 143, 169},
    { 51,  41, 243, 220},
    {219, 116, 223, 251},
    { 18,  26, 216, 218},
    {151,  14,  33, 127},
    { 60,   5, 196, 150},
    {215, 243,  58,  28},
    {174,  63, 157, 118},
    {206, 114,  87,  31},
    {136, 133, 244, 194},
    {186, 229, 173, 213},
    { 41, 179, 177, 144},
    {155, 189,  65, 198},
    { 57, 111, 232, 170},
    { 21, 162, 241,  98},
    {123,  14,  94, 182},
    {187,   8, 254, 152}
  };
  // verilog_format: on

  logic [7:0] msg_reg [64];
  logic       vld_reg;

  logic [7:0] mul     [64] [4];
  logic [7:0] add     [ 4];
  logic [7:0] msg_r2  [64];
  logic [7:0] parity  [ 4];
  logic       valid;

  // Input registers
  always_ff @(posedge clk) begin
    msg_reg <= msg_in;
    vld_reg <= vld_in;
  end

  generate
    for (genvar i = 0; i < 64; i++) begin : g_mul
      for (genvar j = 0; j < 4; j++) begin

        assign mul[i][j] =
          (msg_reg[i][0] ? g_table_a0[i][j] : 8'b0) ^
          (msg_reg[i][1] ? g_table_a1[i][j] : 8'b0) ^
          (msg_reg[i][2] ? g_table_a2[i][j] : 8'b0) ^
          (msg_reg[i][3] ? g_table_a3[i][j] : 8'b0) ^
          (msg_reg[i][4] ? g_table_a4[i][j] : 8'b0) ^
          (msg_reg[i][5] ? g_table_a5[i][j] : 8'b0) ^
          (msg_reg[i][6] ? g_table_a6[i][j] : 8'b0) ^
          (msg_reg[i][7] ? g_table_a7[i][j] : 8'b0);

      end
    end
  endgenerate

  generate
    for (genvar j = 0; j < 4; j++) begin : g_add

      always_comb begin
        add[j] = '0;
        for (int i = 0; i < 64; i++) begin
          add[j] = add[j] ^ mul[i][j];
        end
      end

    end
  endgenerate

  always_ff @(posedge clk) begin
    msg_r2 <= msg_reg;
  end

  assign msg_out = msg_r2;

  generate
    for (genvar j = 0; j < 4; j++) begin : g_parity

      always_ff @(posedge clk) begin
        parity[j] <= add[j];
      end

      assign parity_out[j] = parity[j];

    end
  endgenerate

  always_ff @(posedge clk) begin
    valid <= vld_reg;
  end

  assign vld_out = valid;

endmodule

`default_nettype wire
